ghdl-grt
